module mux2_32b(a,b,s,z);
    input   [31:0] a,b;
    input   s;
    output   [31:0] z;
    
    mux2_1b m0(a[0],b[0],s,z[0]);
    mux2_1b m1(a[1],b[1],s,z[1]);
    mux2_1b m2(a[2],b[2],s,z[2]);
    mux2_1b m3(a[3],b[3],s,z[3]);
    mux2_1b m4(a[4],b[4],s,z[4]);
    mux2_1b m5(a[5],b[5],s,z[5]);
    mux2_1b m6(a[6],b[6],s,z[6]);
    mux2_1b m7(a[7],b[7],s,z[7]);
    mux2_1b m8(a[8],b[8],s,z[8]);
    mux2_1b m9(a[9],b[9],s,z[9]); 
    mux2_1b m10(a[10],b[10],s,z[10]);
    mux2_1b m11(a[11],b[11],s,z[11]);
    mux2_1b m12(a[12],b[12],s,z[12]);
    mux2_1b m13(a[13],b[13],s,z[13]);
    mux2_1b m14(a[14],b[14],s,z[14]);
    mux2_1b m15(a[15],b[15],s,z[15]);
    mux2_1b m16(a[16],b[16],s,z[16]);
    mux2_1b m17(a[17],b[17],s,z[17]);
    mux2_1b m18(a[18],b[18],s,z[18]);
    mux2_1b m19(a[19],b[19],s,z[19]);
    mux2_1b m20(a[20],b[20],s,z[20]);
    mux2_1b m21(a[21],b[21],s,z[21]);
    mux2_1b m22(a[22],b[22],s,z[22]);
    mux2_1b m23(a[23],b[23],s,z[23]);
    mux2_1b m24(a[24],b[24],s,z[24]);
    mux2_1b m25(a[25],b[25],s,z[25]);
    mux2_1b m26(a[26],b[26],s,z[26]);
    mux2_1b m27(a[27],b[27],s,z[27]);
    mux2_1b m28(a[28],b[28],s,z[28]);
    mux2_1b m29(a[29],b[29],s,z[29]);
    mux2_1b m30(a[30],b[30],s,z[30]);
    mux2_1b m31(a[31],b[31],s,z[31]);
endmodule
