module not_1b(a, z);
  input a;
  output z;
  
  assign z = ~a;
endmodule