module and_1b(a, b, z);
  input a, b;
  output z;
  
  assign z = a & b;
endmodule