module ALU_tb;
  reg [31:0] A, B;
  reg [2:0] ALUSEL, COMPSEL;
  reg ADDSEL, ARITHSEL, SIGN;
  wire [31:0] Z;
  wire OVERFLOW, ZERO, CFLAG;
  
  ALU TEST_ALU(
	.a (A),
	.b (B),
	.AddSel (ADDSEL),
	.ArithSel (ARITHSEL),
	.ALUSel (ALUSEL),
	.CompSel (COMPSEL),
	.sign (SIGN),
	.z (Z),
	.overflow (OVERFLOW),
	.zero (ZERO),
	.cflag (CFLAG)
  );
  
  initial begin
	$display("OR TEST\n");
	$monitor("A = %h, B = %h, Z = %h", A, B, Z);
	#0 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b001; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	#5 ADDSEL = 1'b1; ARITHSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 A = 32'h11111111; B = 32'h00000000;
	#5 A = 32'hffffffff; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h11111111;
	#5 A = 32'h11111111; B = 32'h11111111;
	#5 A = 32'hffffffff; B = 32'h11111111;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h11111111; B = 32'hffffffff;
	#5 A = 32'hffffffff; B = 32'hffffffff;
	#5;
	
	$display("\nAND TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b010; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	#5 ADDSEL = 1'b1; ARITHSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 A = 32'h11111111; B = 32'h00000000;
	#5 A = 32'hffffffff; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h11111111;
	#5 A = 32'h11111111; B = 32'h11111111;
	#5 A = 32'hffffffff; B = 32'h11111111;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h11111111; B = 32'hffffffff;
	#5 A = 32'hffffffff; B = 32'hffffffff;
	#5;
	
	$display("\nXOR TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b011; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	#5 ADDSEL = 1'b1; ARITHSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 A = 32'h11111111; B = 32'h00000000;
	#5 A = 32'hffffffff; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h11111111;
	#5 A = 32'h11111111; B = 32'h11111111;
	#5 A = 32'hffffffff; B = 32'h11111111;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h11111111; B = 32'hffffffff;
	#5 A = 32'hffffffff; B = 32'hffffffff;
	#5;
	
	$display("\nLEFT SHIFT TEST\n");
	#5 A = 32'h000000ab; B = 32'h00000000; ALUSEL = 3'b100; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	#5 ADDSEL = 1'b1; ARITHSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 B = 32'h00000001;
	#5 B = 32'h00000011;
	#5 B = 32'h00000110;
	#5 A = 32'h800000ab; B = 32'h00000011;
	#5 A = 32'h80000d2c; B = 32'h00001000;
	#5 B = 32'h00001001;
	#5;
	
	$display("\nRIGHT SHIFT LOGICAL TEST\n");
	#5 A = 32'h000000aa; B = 32'h00000000; ALUSEL = 3'b101; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	#5 ADDSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 B = 32'h00000002;
	#5 A = 32'h00000001; B = 32'h00000003;
	#5 A = 32'h00000011;
	#5 A = 32'h80000000; B = 32'h00000011;
	#5 A = 32'hffff0000; B = 32'h00000005;
	#5;
	$display("\nRIGHT SHIFT ARITHMETIC TEST\n");
	#5 A = 32'h000000aa; B = 32'h00000000; ARITHSEL = 1'b1;
	#5 A = 32'h00000001;
	#5 A = 32'h00000001; B = 32'h00000001;
	#5 A = 32'h00000003;
	#5 A = 32'h80000000; B = 32'h00000005;
	#5 A = 32'hffff0000; B = 32'h00000004;
	#5;
	
	$display("\nUNSIGNED GREATER THAN TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nUNSIGNED GREATER THAN OR EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b001; SIGN = 1'b0;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nUNSIGNED LESS THAN TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b010; SIGN = 1'b0;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nUNSIGNED LESS THAN OR EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b011; SIGN = 1'b0;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nUNSIGNED EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b100; SIGN = 1'b0;
	#5 ARITHSEL = 1'b1; COMPSEL = 3'b110;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nUNSIGNED NOT EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b101; SIGN = 1'b0;
	#5 ARITHSEL = 1'b1; COMPSEL = 3'b111;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nSIGNED GREATER THAN TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b1;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nSIGNED GREATER THAN OR EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b001; SIGN = 1'b1;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nSIGNED LESS THAN TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b010; SIGN = 1'b1;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nSIGNED LESS THAN OR EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b011; SIGN = 1'b1;
	#5 ARITHSEL = 1'b1;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nSIGNED EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b100; SIGN = 1'b1;
	#5 ARITHSEL = 1'b1; COMPSEL = 3'b110;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	$display("\nSIGNED NOT EQUAL TO TEST\n");
	#5 A = 32'h00000000; B = 32'h00000000; ALUSEL = 3'b110; ADDSEL = 1'b1; ARITHSEL = 1'b0; COMPSEL = 3'b101; SIGN = 1'b1;
	#5 ARITHSEL = 1'b1; COMPSEL = 3'b111;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'h0000ffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffff0000;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5 A = 32'h00000000; B = 32'hffffffff;
	#5 A = 32'h0000ffff;
	#5 A = 32'hffff0000;
	#5 A = 32'hffffffff;
	#5;
	
	$display("\nUNSIGNED ADDITION TEST\n");
	$monitor("A = %h, B = %h, Z = %h, CFLAG = %b, ZERO = %b", A, B, Z, CFLAG, ZERO);
	#5 A = 32'h00000014; B = 32'h00000035; ALUSEL = 3'b000; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b0;
	//#5 ARITHSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 A = 32'h00000001; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h00000001;
	#5 A = 32'h00000000; B = 32'h00000000;
	#5 A = 32'h80000000; B = 32'h7fffffff;
	#5 A = 32'h80000000; B = 32'hffffffff;
	#5 A = 32'h00000001; B = 32'hffffffff;
	#5 A = 32'h7fffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h00000001;
	#5 ADDSEL = 1'b1;
	$display("\nUNSIGNED SUBTRACTION TEST\n");
	#5 A = 32'h00000035; B = 32'h00000014; 
	#5 A = 32'h00000010; B = 32'h00000008;
	#5 A = 32'h00000001; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h00000001;
	#5 A = 32'h00000000; B = 32'h00000000;
	#5 A = 32'h80000000; B = 32'h7fffffff;
	#5 A = 32'h80000000; B = 32'hffffffff;
	#5 A = 32'h00000001; B = 32'hffffffff;
	#5 A = 32'h7fffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h00000001;
	#5;

	$display("\nSIGNED ADDITION TEST\n");
	$monitor("A = %h, B = %h, Z = %h, OVERFLOW = %b, ZERO = %b", A, B, Z, OVERFLOW, ZERO);
	#5 A = 32'h00000014; B = 32'h00000035; ALUSEL = 3'b000; ADDSEL = 1'b0; ARITHSEL = 1'b0; COMPSEL = 3'b000; SIGN = 1'b1;
	//#5 ARITHSEL = 1'b1; COMPSEL = 3'b111; SIGN = 1'b1;
	#5 A = 32'h00000001; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h00000001;
	#5 A = 32'h00000000; B = 32'h00000000;
	#5 A = 32'h80000000; B = 32'h7fffffff;
	#5 A = 32'h80000000; B = 32'hffffffff;
	#5 A = 32'h00000001; B = 32'hffffffff;
	#5 A = 32'h7fffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h00000001;
	#5 A = 32'h7fffffff; B = 32'h00000001;
	#5 ADDSEL = 1'b1;
	$display("\nSIGNED SUBTRACTION TEST\n");
	#5 A = 32'h00000035; B = 32'h00000014;
	#5 A = 32'h00000010; B = 32'h00000008;
	#5 A = 32'h00000001; B = 32'h00000000;
	#5 A = 32'h00000000; B = 32'h00000001;
	#5 A = 32'h00000000; B = 32'h00000000;
	#5 A = 32'h80000000; B = 32'h7fffffff;
	#5 A = 32'h80000000; B = 32'hffffffff;
	#5 A = 32'h00000001; B = 32'hffffffff;
	#5 A = 32'h7fffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h80000000;
	#5 A = 32'hffffffff; B = 32'h00000001;
	#5;
  end
endmodule
