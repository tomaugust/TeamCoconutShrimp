module mux8_32b_tb;
    reg [31:0] A;
    reg [31:0] B;
    reg [31:0] C;
    reg [31:0] D;
    reg [31:0] E;
    reg [31:0] F;
    reg [31:0] G;
    reg [31:0] H;
    reg [2:0]SEL;
    wire [31:0] Z;
    
    mux8_32b MUX8_32B(.a(A),.b(B),.c(C),.d(D),.e(E),.f(F),.g(G),.h(H),.s(SEL),.z(Z));
    
    initial begin
        $monitor("A=%h B=%h C=%h D=%h E=%h F=%h G=%h H=%h SEL=%b Z=%h",A,B,C,D,E,F,G,H,SEL,Z);
        #0 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444 ;F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b000;
        #1 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b001;
        #1 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b010;
        #1 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b011;
        #1 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b100;
        #1 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b101;
        #1 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b110;
        #2 A=32'h00000000; B=32'h11111111; C=32'h22222222; D=32'h33333333; E=32'h44444444; F=32'h55555555; G=32'h66666666; H=32'h77777777; SEL=3'b111;
    end
endmodule
